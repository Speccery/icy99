// tms9918_tb.v
`timescale 1ns / 1ns

module tms9918_tb();

reg clk=1'b0, reset=1'b1, 
    mode=1'b0;  // 1=reg 0=memory
reg [7:0] vdp_addr;
reg [7:0] vdp_data_in;
wire [15:0] vdp_data_out;
reg wr=1'b0;
reg rd=1'b0;
wire vga_vsync, vga_hsync;
wire debug1, debug2, int_out;
wire [2:0] vga_red, vga_green;
wire [1:0] vga_blue;

tms9918 DUT(
    .clk(clk),
    .reset(reset),
    .mode(mode),
    .addr(vdp_addr),
    .data_in(vdp_data_in),
    .data_out(vdp_data_out),
    .wr(wr),
    .rd(rd),
    .vga_vsync(vga_vsync),
    .vga_hsync(vga_hsync),
    .debug1(debug1),
    .debug2(debug2),
    .int_out(int_out),
    .vga_red(vga_red),
    .vga_green(vga_green),
    .vga_blue(vga_blue)
);

// 25MHz clock, 40 ns cycle time, toggle every half cycle
always #20 clk = !clk;   

reg [7:0] my_count = 0;

initial begin
    // EP testing location of vcd file - put it to /tmp so it does not get synced by Dropbox
    $dumpfile("sim-tms9918_tb.lxt"); // iverilog -lxt2 argument
//    $dumpfile("/tmp/tms9918_tb.vcd");
    $dumpvars(0, tms9918_tb);
    $display("tms9918_tb started");
    #500 reset = 1'b0;
    #500

    // Initialize the VDP
    vdp_init();

    // Write one font description to 0x800
    mode = 1;
    vdp_write(0, 8'h00);
    vdp_write(0, 8'h40 | 8'h08);    // Setup write to 0x0800
    @(posedge clk)
      ;
    mode = 0;
    vdp_write(0, 8'b0000_0000); // write the actual data
    vdp_write(0, 8'b0111_0000); 
    vdp_write(0, 8'b1000_1000); 
    vdp_write(0, 8'b1111_1000);
    vdp_write(0, 8'b1000_1000); 
    vdp_write(0, 8'b1000_1000);
    vdp_write(0, 8'b1000_1000); 
    vdp_write(0, 8'b1000_1000);

    // Write the first row of characters
    mode = 1;
    vdp_write(0, 8'h00);
    vdp_write(0, 8'h40 | 8'h00);    // Setup write to 0x0000

    mode = 0;
    write_zeros(80);  // write 80 zero bytes.

    mode = 1;
    vdp_write(0, 8'h34);
    vdp_write(0, 8'h40 | 8'h12);    // Setup write to 0x1234
    mode = 0;
    vdp_write(0, 8'h5a); // write the actual data
    vdp_write(0, 8'hee);    // write second databyte
    #100
    // prepare to read back the data
    mode = 1;
    vdp_write(0, 8'h34);
    vdp_write(0, 8'h00 | 8'h12);    // Setup read from 0x1234
    mode = 0;

    #50 rd = 1'b1;
    #150 $display("data read %x\n", vdp_data_out);
    rd = 1'b0;

    #50 rd = 1'b1;
    #150 $display("data read %x\n", vdp_data_out);
    rd = 1'b0;

    #50
    // #100000
    #20000000

    $finish;
end


  task vdp_write;
    input [7:0] waddr;
    input [7:0] wdata;
  
    begin 
        wr = 1'b0;
        vdp_data_in = wdata;
        vdp_addr = waddr;
        @(negedge clk)
          ;
        wr = 1'b1;
        @(posedge clk)
          ;
        wr = 1'b0;
        #50;
    end
  endtask

  task write_zeros;
    input[7:0] count;
    reg[7:0] i;
    begin
      for(i=0; i<count; i++)
        vdp_write(0,0);
    end
  endtask

  task vdp_init;
    begin
      mode = 1;  // Basically the address input, register access
/*
      // Init as TurboForth, 40 column text mode.
      vdp_write(0, 8'h00);    vdp_write(0, 8'h80);  // Reg 0
      vdp_write(0, 8'hF0);    vdp_write(0, 8'h81);  // Reg 1
      vdp_write(0, 8'h00);    vdp_write(0, 8'h82);  // Reg 2
      vdp_write(0, 8'h0E);    vdp_write(0, 8'h83);  // Reg 3
      vdp_write(0, 8'h01);    vdp_write(0, 8'h84);  // Reg 4
      vdp_write(0, 8'h06);    vdp_write(0, 8'h85);  // Reg 5
      vdp_write(0, 8'h00);    vdp_write(0, 8'h86);  // Reg 6
      vdp_write(0, 8'hF4);    vdp_write(0, 8'h87);  // Reg 7
*/    

      // Init as in TI Invaders
      // regs= [ 0x00, 0xE2, 0xF0, 0x0E, 0xF9, 0x86, 0xF8, 0xF1 ]
      vdp_write(0, 8'h00);    vdp_write(0, 8'h80);  // Reg 0
      vdp_write(0, 8'hE2);    vdp_write(0, 8'h81);  // Reg 1
      vdp_write(0, 8'hF0);    vdp_write(0, 8'h82);  // Reg 2
      vdp_write(0, 8'h0E);    vdp_write(0, 8'h83);  // Reg 3
      vdp_write(0, 8'hF9);    vdp_write(0, 8'h84);  // Reg 4
      vdp_write(0, 8'h86);    vdp_write(0, 8'h85);  // Reg 5
      vdp_write(0, 8'hF8);    vdp_write(0, 8'h86);  // Reg 6
      // Changed to F2 to have a different color for border than black
      vdp_write(0, 8'hF2);    vdp_write(0, 8'h87);  // Reg 7

    end
  endtask

endmodule
